`define PDU_IMEM_FILE "your_path_to_pdu_inits/pdu_imem.ini"
`define PDU_DMEM_FILE "your_path_to_pdu_inits/pdu_dmem.ini"
`define CPU_IMEM_FILE "your_path_to_cpu_inits/instr.ini"
`define CPU_DMEM_FILE "your_path_to_cpu_inits/data.ini"